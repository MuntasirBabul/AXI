`ifndef PROJECT_UVM_DEFINES
`define PROJECT_UVM_DEFINES


`endif
